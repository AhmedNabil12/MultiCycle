--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   22:30:51 06/09/2021
-- Design Name:   
-- Module Name:   D:/Computer Arche Lab/ProjectWeek1/MIPSSingleCycle.vhd
-- Project Name:  ProjectWeek1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: MIPS
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY MIPSSingleCycle IS
END MIPSSingleCycle;
 
ARCHITECTURE behavior OF MIPSSingleCycle IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
  COMPONENT MIPS
    PORT(
         reset : IN  std_logic;
         clk : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal reset : std_logic := '0';
   signal clk  COMPONENT MIPS
    PORT(
         reset : IN  std_logic;
         clk_Main : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal reset : std_logic := '0';
   signal clk_Main : std_logic := '0';

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: MIPS PORT MAP (
          reset => reset,
          clk => clk_Main
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk_Main <= '0';
		wait for clk_period/2;
		clk_Main <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
 : std_logic := '0';

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: MIPS PORT MAP (
          reset => reset,
          clk_Main => clk_Main
        );

   -- Clock process definitions
   clk_Main_process :process
   begin
		clk_Main <= '0';
		wait for clk_Main_period/2;
		clk_Main <= '1';
		wait for clk_Main_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_Main_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
